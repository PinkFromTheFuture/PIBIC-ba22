--------------------------------------------------------------
-- ROM_ba22 - Template
-- Author: Renato Sampaio
-- Date: 21/02/2013
--------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;		 
use ieee.std_logic_unsigned.all;

entity ROM_ba22 is
generic(
	ADDR_WIDTH : integer := 14
);
port(	clk   : in std_logic;
		addr	: in std_logic_vector(ADDR_WIDTH-1 downto 0);
		data_out: out std_logic_vector(31 downto 0)
);
end ROM_ba22;

--------------------------------------------------------------

architecture Behav of ROM_ba22 is

    type ROM_Array is array (0 to (2**ADDR_WIDTH)-1 ) 
	of std_logic_vector(31 downto 0);

    constant dados: ROM_Array := (
		0 => "00000000000000000000000000000000",
		1 => "00000000000000000000000000000000",
		2 => "00000000000000000000000000000000",
		3 => "00000000000000000000000000000000",
		4 => "00000000000000000000000000000000",
		5 => "00000000000000000000000000000000",
		6 => "00000000000000000000000000000000",
		7 => "00000000000000000000000000000000",
		8 => "00000000000000000000000000000000",
		9 => "00000000000000000000000000000000",
		10 => "00000000000000000000000000000000",
		11 => "00000000000000000000000000000000",
		12 => "00000000000000000000000000000000",
		13 => "00000000000000000000000000000000",
		14 => "00000000000000000000000000000000",
		15 => "00000000000000000000000000000000",
		16 => "00000000000000000000000000000000",
		17 => "00000000000000000000000000000000",
		18 => "00000000000000000000000000000000",
		19 => "00000000000000000000000000000000",
		20 => "00000000000000000000000000000000",
		21 => "00000000000000000000000000000000",
		22 => "00000000000000000000000000000000",
		23 => "00000000000000000000000000000000",
		24 => "00000000000000000000000000000000",
		25 => "00000000000000000000000000000000",
		26 => "00000000000000000000000000000000",
		27 => "00000000000000000000000000000000",
		28 => "00000000000000000000000000000000",
		29 => "00000000000000000000000000000000",
		30 => "00000000000000000000000000000000",
		31 => "00000000000000000000000000000000",
		32 => "00000000000000000000000000000000",
		33 => "00000000000000000000000000000000",
		34 => "00000000000000000000000000000000",
		35 => "00000000000000000000000000000000",
		36 => "00000000000000000000000000000000",
		37 => "00000000000000000000000000000000",
		38 => "00000000000000000000000000000000",
		39 => "00000000000000000000000000000000",
		40 => "00000000000000000000000000000000",
		41 => "00000000000000000000000000000000",
		42 => "00000000000000000000000000000000",
		43 => "00000000000000000000000000000000",
		44 => "00000000000000000000000000000000",
		45 => "00000000000000000000000000000000",
		46 => "00000000000000000000000000000000",
		47 => "00000000000000000000000000000000",
		48 => "00000000000000000000000000000000",
		49 => "00000000000000000000000000000000",
		50 => "00000000000000000000000000000000",
		51 => "00000000000000000000000000000000",
		52 => "00000000000000000000000000000000",
		53 => "00000000000000000000000000000000",
		54 => "00000000000000000000000000000000",
		55 => "00000000000000000000000000000000",
		56 => "00000000000000000000000000000000",
		57 => "00000000000000000000000000000000",
		58 => "00000000000000000000000000000000",
		59 => "00000000000000000000000000000000",
		60 => "00000000000000000000000000000000",
		61 => "00000000000000000000000000000000",
		62 => "00000000000000000000000000000000",
		63 => "00000000000000000000000000000000",
		64 => "10011000001000000011111111111100",
		65 => "00000000000000001001010000100001",
		66 => "00011111111111111111111111111111",
		67 => "10011000011000000010001100000100",
		68 => "00000000000000001001100010000000",
		69 => "00100011000001000000000000000000",
		70 => "01001011111000000000000010011000",
		71 => "01100000001011010000010000000000",
		72 => "00000000100110001000000000101101",
		73 => "00000100000000000000000001001000",
		74 => "00100000000000001001100001000000",
		75 => "00101101000001010000000000000000",
		76 => "01001000011111011110000000000000",
		77 => "00011000000011011111111111010011",
		78 => "10000110010010111000000000000000",
		79 => "01110010110100111100011001000101",
		80 => "00000000110011000000001100111111",
		81 => "11111111000011011011111100000000",
		82 => "01110011110100111000011001001101",
		83 => "00000000001000000000001100000000",
		84 => "00000000011110000000111110111111",
		85 => "01000111110100000000000000000000",
		86 => "00000000000000000000000000000000",
		87 => "00000000000000000000000000000000",
		88 => "00000000000000000000000000000000",
		89 => "00000000000000000000000000000000",
		90 => "00000000000000000000000000000000",
		91 => "00000000000000000000000000000000",
		92 => "00000000000000000000000000000000",
		93 => "00000000000000000000000000000000",
		94 => "00000000000000000000000000000000",
		95 => "00000000000000000000000000000000",
		96 => "00000000000000000000000000000000",
		97 => "00000000000000000000000000000000",
		98 => "00000000000000000000000000000000",
		99 => "00000000000000000000000000000000",
		100 => "00000000000000000000000000000000",
		101 => "00000000000000000000000000000000",
		102 => "00000000000000000000000000000000",
		103 => "00000000000000000000000000000000",
		104 => "00000000000000000000000000000000",
		105 => "00000000000000000000000000000000",
		106 => "00000000000000000000000000000000",
		107 => "00000000000000000000000000000000",
		108 => "00000000000000000000000000000000",
		109 => "00000000000000000000000000000000",
		110 => "00000000000000000000000000000000",
		111 => "00000000000000000000000000000000",
		112 => "00000000000000000000000000000000",
		113 => "00000000000000000000000000000000",
		114 => "00000000000000000000000000000000",
		115 => "00000000000000000000000000000000",
		116 => "00000000000000000000000000000000",
		117 => "00000000000000000000000000000000",
		118 => "00000000000000000000000000000000",
		119 => "00000000000000000000000000000000",
		120 => "00000000000000000000000000000000",
		121 => "00000000000000000000000000000000",
		122 => "00000000000000000000000000000000",
		123 => "00000000000000000000000000000000",
		124 => "00000000000000000000000000000000",
		125 => "00000000000000000000000000000000",
		126 => "00000000000000000000000000000000",
		127 => "00000000000000000000000000000000",
		128 => "00000000000110000000010000000000",
		129 => "00000000000000000000000000000000",
		130 => "00000000000000000000000000000000",
		131 => "00000000000000000000000000000000",
		132 => "00000000000000000000000000000000",
		133 => "00000000000000000000000000000000",
		134 => "00000000000000000000000000000000",
		135 => "00000000000000000000000000000000",
		136 => "00000000000000000000000000000000",
		137 => "00000000000000000000000000000000",
		138 => "00000000000000000000000000000000",
		139 => "00000000000000000000000000000000",
		140 => "00000000000000000000000000000000",
		141 => "00000000000000000000000000000000",
		142 => "00000000000000000000000000000000",
		143 => "00000000000000000000000000000000",
		144 => "00000000000000000000000000000000",
		145 => "00000000000000000000000000000000",
		146 => "00000000000000000000000000000000",
		147 => "00000000000000000000000000000000",
		148 => "00000000000000000000000000000000",
		149 => "00000000000000000000000000000000",
		150 => "00000000000000000000000000000000",
		151 => "00000000000000000000000000000000",
		152 => "00000000000000000000000000000000",
		153 => "00000000000000000000000000000000",
		154 => "00000000000000000000000000000000",
		155 => "00000000000000000000000000000000",
		156 => "00000000000000000000000000000000",
		157 => "00000000000000000000000000000000",
		158 => "00000000000000000000000000000000",
		159 => "00000000000000000000000000000000",
		160 => "00000000000000000000000000000000",
		161 => "00000000000000000000000000000000",
		162 => "00000000000000000000000000000000",
		163 => "00000000000000000000000000000000",
		164 => "00000000000000000000000000000000",
		165 => "00000000000000000000000000000000",
		166 => "00000000000000000000000000000000",
		167 => "00000000000000000000000000000000",
		168 => "00000000000000000000000000000000",
		169 => "00000000000000000000000000000000",
		170 => "00000000000000000000000000000000",
		171 => "00000000000000000000000000000000",
		172 => "00000000000000000000000000000000",
		173 => "00000000000000000000000000000000",
		174 => "00000000000000000000000000000000",
		175 => "00000000000000000000000000000000",
		176 => "00000000000000000000000000000000",
		177 => "00000000000000000000000000000000",
		178 => "00000000000000000000000000000000",
		179 => "00000000000000000000000000000000",
		180 => "00000000000000000000000000000000",
		181 => "00000000000000000000000000000000",
		182 => "00000000000000000000000000000000",
		183 => "00000000000000000000000000000000",
		184 => "00000000000000000000000000000000",
		185 => "00000000000000000000000000000000",
		186 => "00000000000000000000000000000000",
		187 => "00000000000000000000000000000000",
		188 => "00000000000000000000000000000000",
		189 => "00000000000000000000000000000000",
		190 => "00000000000000000000000000000000",
		191 => "00000000000000000000000000000000",
		192 => "00000000000110000000010000000000",
		193 => "00000000000000000000000000000000",
		194 => "00000000000000000000000000000000",
		195 => "00000000000000000000000000000000",
		196 => "00000000000000000000000000000000",
		197 => "00000000000000000000000000000000",
		198 => "00000000000000000000000000000000",
		199 => "00000000000000000000000000000000",
		200 => "00000000000000000000000000000000",
		201 => "00000000000000000000000000000000",
		202 => "00000000000000000000000000000000",
		203 => "00000000000000000000000000000000",
		204 => "00000000000000000000000000000000",
		205 => "00000000000000000000000000000000",
		206 => "00000000000000000000000000000000",
		207 => "00000000000000000000000000000000",
		208 => "00000000000000000000000000000000",
		209 => "00000000000000000000000000000000",
		210 => "00000000000000000000000000000000",
		211 => "00000000000000000000000000000000",
		212 => "00000000000000000000000000000000",
		213 => "00000000000000000000000000000000",
		214 => "00000000000000000000000000000000",
		215 => "00000000000000000000000000000000",
		216 => "00000000000000000000000000000000",
		217 => "00000000000000000000000000000000",
		218 => "00000000000000000000000000000000",
		219 => "00000000000000000000000000000000",
		220 => "00000000000000000000000000000000",
		221 => "00000000000000000000000000000000",
		222 => "00000000000000000000000000000000",
		223 => "00000000000000000000000000000000",
		224 => "00000000000000000000000000000000",
		225 => "00000000000000000000000000000000",
		226 => "00000000000000000000000000000000",
		227 => "00000000000000000000000000000000",
		228 => "00000000000000000000000000000000",
		229 => "00000000000000000000000000000000",
		230 => "00000000000000000000000000000000",
		231 => "00000000000000000000000000000000",
		232 => "00000000000000000000000000000000",
		233 => "00000000000000000000000000000000",
		234 => "00000000000000000000000000000000",
		235 => "00000000000000000000000000000000",
		236 => "00000000000000000000000000000000",
		237 => "00000000000000000000000000000000",
		238 => "00000000000000000000000000000000",
		239 => "00000000000000000000000000000000",
		240 => "00000000000000000000000000000000",
		241 => "00000000000000000000000000000000",
		242 => "00000000000000000000000000000000",
		243 => "00000000000000000000000000000000",
		244 => "00000000000000000000000000000000",
		245 => "00000000000000000000000000000000",
		246 => "00000000000000000000000000000000",
		247 => "00000000000000000000000000000000",
		248 => "00000000000000000000000000000000",
		249 => "00000000000000000000000000000000",
		250 => "00000000000000000000000000000000",
		251 => "00000000000000000000000000000000",
		252 => "00000000000000000000000000000000",
		253 => "00000000000000000000000000000000",
		254 => "00000000000000000000000000000000",
		255 => "00000000000000000000000000000000",
		256 => "00000000000110000000010000000000",
		257 => "00000000000000000000000000000000",
		258 => "00000000000000000000000000000000",
		259 => "00000000000000000000000000000000",
		260 => "00000000000000000000000000000000",
		261 => "00000000000000000000000000000000",
		262 => "00000000000000000000000000000000",
		263 => "00000000000000000000000000000000",
		264 => "00000000000000000000000000000000",
		265 => "00000000000000000000000000000000",
		266 => "00000000000000000000000000000000",
		267 => "00000000000000000000000000000000",
		268 => "00000000000000000000000000000000",
		269 => "00000000000000000000000000000000",
		270 => "00000000000000000000000000000000",
		271 => "00000000000000000000000000000000",
		272 => "00000000000000000000000000000000",
		273 => "00000000000000000000000000000000",
		274 => "00000000000000000000000000000000",
		275 => "00000000000000000000000000000000",
		276 => "00000000000000000000000000000000",
		277 => "00000000000000000000000000000000",
		278 => "00000000000000000000000000000000",
		279 => "00000000000000000000000000000000",
		280 => "00000000000000000000000000000000",
		281 => "00000000000000000000000000000000",
		282 => "00000000000000000000000000000000",
		283 => "00000000000000000000000000000000",
		284 => "00000000000000000000000000000000",
		285 => "00000000000000000000000000000000",
		286 => "00000000000000000000000000000000",
		287 => "00000000000000000000000000000000",
		288 => "00000000000000000000000000000000",
		289 => "00000000000000000000000000000000",
		290 => "00000000000000000000000000000000",
		291 => "00000000000000000000000000000000",
		292 => "00000000000000000000000000000000",
		293 => "00000000000000000000000000000000",
		294 => "00000000000000000000000000000000",
		295 => "00000000000000000000000000000000",
		296 => "00000000000000000000000000000000",
		297 => "00000000000000000000000000000000",
		298 => "00000000000000000000000000000000",
		299 => "00000000000000000000000000000000",
		300 => "00000000000000000000000000000000",
		301 => "00000000000000000000000000000000",
		302 => "00000000000000000000000000000000",
		303 => "00000000000000000000000000000000",
		304 => "00000000000000000000000000000000",
		305 => "00000000000000000000000000000000",
		306 => "00000000000000000000000000000000",
		307 => "00000000000000000000000000000000",
		308 => "00000000000000000000000000000000",
		309 => "00000000000000000000000000000000",
		310 => "00000000000000000000000000000000",
		311 => "00000000000000000000000000000000",
		312 => "00000000000000000000000000000000",
		313 => "00000000000000000000000000000000",
		314 => "00000000000000000000000000000000",
		315 => "00000000000000000000000000000000",
		316 => "00000000000000000000000000000000",
		317 => "00000000000000000000000000000000",
		318 => "00000000000000000000000000000000",
		319 => "00000000000000000000000000000000",
		320 => "00000000000110000000010000000000",
		321 => "00000000000000000000000000000000",
		322 => "00000000000000000000000000000000",
		323 => "00000000000000000000000000000000",
		324 => "00000000000000000000000000000000",
		325 => "00000000000000000000000000000000",
		326 => "00000000000000000000000000000000",
		327 => "00000000000000000000000000000000",
		328 => "00000000000000000000000000000000",
		329 => "00000000000000000000000000000000",
		330 => "00000000000000000000000000000000",
		331 => "00000000000000000000000000000000",
		332 => "00000000000000000000000000000000",
		333 => "00000000000000000000000000000000",
		334 => "00000000000000000000000000000000",
		335 => "00000000000000000000000000000000",
		336 => "00000000000000000000000000000000",
		337 => "00000000000000000000000000000000",
		338 => "00000000000000000000000000000000",
		339 => "00000000000000000000000000000000",
		340 => "00000000000000000000000000000000",
		341 => "00000000000000000000000000000000",
		342 => "00000000000000000000000000000000",
		343 => "00000000000000000000000000000000",
		344 => "00000000000000000000000000000000",
		345 => "00000000000000000000000000000000",
		346 => "00000000000000000000000000000000",
		347 => "00000000000000000000000000000000",
		348 => "00000000000000000000000000000000",
		349 => "00000000000000000000000000000000",
		350 => "00000000000000000000000000000000",
		351 => "00000000000000000000000000000000",
		352 => "00000000000000000000000000000000",
		353 => "00000000000000000000000000000000",
		354 => "00000000000000000000000000000000",
		355 => "00000000000000000000000000000000",
		356 => "00000000000000000000000000000000",
		357 => "00000000000000000000000000000000",
		358 => "00000000000000000000000000000000",
		359 => "00000000000000000000000000000000",
		360 => "00000000000000000000000000000000",
		361 => "00000000000000000000000000000000",
		362 => "00000000000000000000000000000000",
		363 => "00000000000000000000000000000000",
		364 => "00000000000000000000000000000000",
		365 => "00000000000000000000000000000000",
		366 => "00000000000000000000000000000000",
		367 => "00000000000000000000000000000000",
		368 => "00000000000000000000000000000000",
		369 => "00000000000000000000000000000000",
		370 => "00000000000000000000000000000000",
		371 => "00000000000000000000000000000000",
		372 => "00000000000000000000000000000000",
		373 => "00000000000000000000000000000000",
		374 => "00000000000000000000000000000000",
		375 => "00000000000000000000000000000000",
		376 => "00000000000000000000000000000000",
		377 => "00000000000000000000000000000000",
		378 => "00000000000000000000000000000000",
		379 => "00000000000000000000000000000000",
		380 => "00000000000000000000000000000000",
		381 => "00000000000000000000000000000000",
		382 => "00000000000000000000000000000000",
		383 => "00000000000000000000000000000000",
		384 => "00000000000110000000010000000000",
		385 => "00000000000000000000000000000000",
		386 => "00000000000000000000000000000000",
		387 => "00000000000000000000000000000000",
		388 => "00000000000000000000000000000000",
		389 => "00000000000000000000000000000000",
		390 => "00000000000000000000000000000000",
		391 => "00000000000000000000000000000000",
		392 => "00000000000000000000000000000000",
		393 => "00000000000000000000000000000000",
		394 => "00000000000000000000000000000000",
		395 => "00000000000000000000000000000000",
		396 => "00000000000000000000000000000000",
		397 => "00000000000000000000000000000000",
		398 => "00000000000000000000000000000000",
		399 => "00000000000000000000000000000000",
		400 => "00000000000000000000000000000000",
		401 => "00000000000000000000000000000000",
		402 => "00000000000000000000000000000000",
		403 => "00000000000000000000000000000000",
		404 => "00000000000000000000000000000000",
		405 => "00000000000000000000000000000000",
		406 => "00000000000000000000000000000000",
		407 => "00000000000000000000000000000000",
		408 => "00000000000000000000000000000000",
		409 => "00000000000000000000000000000000",
		410 => "00000000000000000000000000000000",
		411 => "00000000000000000000000000000000",
		412 => "00000000000000000000000000000000",
		413 => "00000000000000000000000000000000",
		414 => "00000000000000000000000000000000",
		415 => "00000000000000000000000000000000",
		416 => "00000000000000000000000000000000",
		417 => "00000000000000000000000000000000",
		418 => "00000000000000000000000000000000",
		419 => "00000000000000000000000000000000",
		420 => "00000000000000000000000000000000",
		421 => "00000000000000000000000000000000",
		422 => "00000000000000000000000000000000",
		423 => "00000000000000000000000000000000",
		424 => "00000000000000000000000000000000",
		425 => "00000000000000000000000000000000",
		426 => "00000000000000000000000000000000",
		427 => "00000000000000000000000000000000",
		428 => "00000000000000000000000000000000",
		429 => "00000000000000000000000000000000",
		430 => "00000000000000000000000000000000",
		431 => "00000000000000000000000000000000",
		432 => "00000000000000000000000000000000",
		433 => "00000000000000000000000000000000",
		434 => "00000000000000000000000000000000",
		435 => "00000000000000000000000000000000",
		436 => "00000000000000000000000000000000",
		437 => "00000000000000000000000000000000",
		438 => "00000000000000000000000000000000",
		439 => "00000000000000000000000000000000",
		440 => "00000000000000000000000000000000",
		441 => "00000000000000000000000000000000",
		442 => "00000000000000000000000000000000",
		443 => "00000000000000000000000000000000",
		444 => "00000000000000000000000000000000",
		445 => "00000000000000000000000000000000",
		446 => "00000000000000000000000000000000",
		447 => "00000000000000000000000000000000",
		448 => "00000000000110000000010000000000",
		449 => "00000000000000000000000000000000",
		450 => "00000000000000000000000000000000",
		451 => "00000000000000000000000000000000",
		452 => "00000000000000000000000000000000",
		453 => "00000000000000000000000000000000",
		454 => "00000000000000000000000000000000",
		455 => "00000000000000000000000000000000",
		456 => "00000000000000000000000000000000",
		457 => "00000000000000000000000000000000",
		458 => "00000000000000000000000000000000",
		459 => "00000000000000000000000000000000",
		460 => "00000000000000000000000000000000",
		461 => "00000000000000000000000000000000",
		462 => "00000000000000000000000000000000",
		463 => "00000000000000000000000000000000",
		464 => "00000000000000000000000000000000",
		465 => "00000000000000000000000000000000",
		466 => "00000000000000000000000000000000",
		467 => "00000000000000000000000000000000",
		468 => "00000000000000000000000000000000",
		469 => "00000000000000000000000000000000",
		470 => "00000000000000000000000000000000",
		471 => "00000000000000000000000000000000",
		472 => "00000000000000000000000000000000",
		473 => "00000000000000000000000000000000",
		474 => "00000000000000000000000000000000",
		475 => "00000000000000000000000000000000",
		476 => "00000000000000000000000000000000",
		477 => "00000000000000000000000000000000",
		478 => "00000000000000000000000000000000",
		479 => "00000000000000000000000000000000",
		480 => "00000000000000000000000000000000",
		481 => "00000000000000000000000000000000",
		482 => "00000000000000000000000000000000",
		483 => "00000000000000000000000000000000",
		484 => "00000000000000000000000000000000",
		485 => "00000000000000000000000000000000",
		486 => "00000000000000000000000000000000",
		487 => "00000000000000000000000000000000",
		488 => "00000000000000000000000000000000",
		489 => "00000000000000000000000000000000",
		490 => "00000000000000000000000000000000",
		491 => "00000000000000000000000000000000",
		492 => "00000000000000000000000000000000",
		493 => "00000000000000000000000000000000",
		494 => "00000000000000000000000000000000",
		495 => "00000000000000000000000000000000",
		496 => "00000000000000000000000000000000",
		497 => "00000000000000000000000000000000",
		498 => "00000000000000000000000000000000",
		499 => "00000000000000000000000000000000",
		500 => "00000000000000000000000000000000",
		501 => "00000000000000000000000000000000",
		502 => "00000000000000000000000000000000",
		503 => "00000000000000000000000000000000",
		504 => "00000000000000000000000000000000",
		505 => "00000000000000000000000000000000",
		506 => "00000000000000000000000000000000",
		507 => "00000000000000000000000000000000",
		508 => "00000000000000000000000000000000",
		509 => "00000000000000000000000000000000",
		510 => "00000000000000000000000000000000",
		511 => "00000000000000000000000000000000",
		512 => "11001100001000010001110011111111",
		513 => "11011000001000010001110011111111",
		514 => "01010100010000011010000001010100",
		515 => "10100001100010000101010100000001",
		516 => "11111000101010011010000000000100",
		517 => "00000000000000000000000010101001",
		518 => "11000000000000100000000000000000",
		519 => "00000000101010011110000000001100",
		520 => "00000000000000000000000001010101",
		521 => "10100001101111000000010001100001",
		522 => "01001000011011111010000001010001",
		523 => "10100001101111001010100110100000",
		524 => "00000100000000000000000000000001",
		525 => "10101001110000000000001000000000",
		526 => "00000000000000011010100111100000",
		527 => "00001100000000000000000000000001",
		528 => "01010000010000011010000001010000",
		529 => "10100001100010000101000100000001",
		530 => "11111000001011000010000101000000",
		531 => "00000100000000000000000000000000",
		532 => "00000000000000000000000000000000",
		533 => "00000000000000000000000000000000",
		534 => "00000000000000000000000000000000",
		535 => "00000000000000000000000000000000",
		536 => "00000000000000000000000000000000",
		537 => "00000000000000000000000000000000",
		538 => "00000000000000000000000000000000",
		539 => "00000000000000000000000000000000",
		540 => "00000000000000000000000000000000",
		541 => "00000000000000000000000000000000",
		542 => "00000000000000000000000000000000",
		543 => "00000000000000000000000000000000",
		544 => "00000000000000000000000000000000",
		545 => "00000000000000000000000000000000",
		546 => "00000000000000000000000000000000",
		547 => "00000000000000000000000000000000",
		548 => "00000000000000000000000000000000",
		549 => "00000000000000000000000000000000",
		550 => "00000000000000000000000000000000",
		551 => "00000000000000000000000000000000",
		552 => "00000000000000000000000000000000",
		553 => "00000000000000000000000000000000",
		554 => "00000000000000000000000000000000",
		555 => "00000000000000000000000000000000",
		556 => "00000000000000000000000000000000",
		557 => "00000000000000000000000000000000",
		558 => "00000000000000000000000000000000",
		559 => "00000000000000000000000000000000",
		560 => "00000000000000000000000000000000",
		561 => "00000000000000000000000000000000",
		562 => "00000000000000000000000000000000",
		563 => "00000000000000000000000000000000",
		564 => "00000000000000000000000000000000",
		565 => "00000000000000000000000000000000",
		566 => "00000000000000000000000000000000",
		567 => "00000000000000000000000000000000",
		568 => "00000000000000000000000000000000",
		569 => "00000000000000000000000000000000",
		570 => "00000000000000000000000000000000",
		571 => "00000000000000000000000000000000",
		572 => "00000000000000000000000000000000",
		573 => "00000000000000000000000000000000",
		574 => "00000000000000000000000000000000",
		575 => "00000000000000000000000000000000",
		576 => "00000000000110000000010000000000",
		577 => "00000000000000000000000000000000",
		578 => "00000000000000000000000000000000",
		579 => "00000000000000000000000000000000",
		580 => "00000000000000000000000000000000",
		581 => "00000000000000000000000000000000",
		582 => "00000000000000000000000000000000",
		583 => "00000000000000000000000000000000",
		584 => "00000000000000000000000000000000",
		585 => "00000000000000000000000000000000",
		586 => "00000000000000000000000000000000",
		587 => "00000000000000000000000000000000",
		588 => "00000000000000000000000000000000",
		589 => "00000000000000000000000000000000",
		590 => "00000000000000000000000000000000",
		591 => "00000000000000000000000000000000",
		592 => "00000000000000000000000000000000",
		593 => "00000000000000000000000000000000",
		594 => "00000000000000000000000000000000",
		595 => "00000000000000000000000000000000",
		596 => "00000000000000000000000000000000",
		597 => "00000000000000000000000000000000",
		598 => "00000000000000000000000000000000",
		599 => "00000000000000000000000000000000",
		600 => "00000000000000000000000000000000",
		601 => "00000000000000000000000000000000",
		602 => "00000000000000000000000000000000",
		603 => "00000000000000000000000000000000",
		604 => "00000000000000000000000000000000",
		605 => "00000000000000000000000000000000",
		606 => "00000000000000000000000000000000",
		607 => "00000000000000000000000000000000",
		608 => "00000000000000000000000000000000",
		609 => "00000000000000000000000000000000",
		610 => "00000000000000000000000000000000",
		611 => "00000000000000000000000000000000",
		612 => "00000000000000000000000000000000",
		613 => "00000000000000000000000000000000",
		614 => "00000000000000000000000000000000",
		615 => "00000000000000000000000000000000",
		616 => "00000000000000000000000000000000",
		617 => "00000000000000000000000000000000",
		618 => "00000000000000000000000000000000",
		619 => "00000000000000000000000000000000",
		620 => "00000000000000000000000000000000",
		621 => "00000000000000000000000000000000",
		622 => "00000000000000000000000000000000",
		623 => "00000000000000000000000000000000",
		624 => "00000000000000000000000000000000",
		625 => "00000000000000000000000000000000",
		626 => "00000000000000000000000000000000",
		627 => "00000000000000000000000000000000",
		628 => "00000000000000000000000000000000",
		629 => "00000000000000000000000000000000",
		630 => "00000000000000000000000000000000",
		631 => "00000000000000000000000000000000",
		632 => "00000000000000000000000000000000",
		633 => "00000000000000000000000000000000",
		634 => "00000000000000000000000000000000",
		635 => "00000000000000000000000000000000",
		636 => "00000000000000000000000000000000",
		637 => "00000000000000000000000000000000",
		638 => "00000000000000000000000000000000",
		639 => "00000000000000000000000000000000",
		640 => "00000000000110000000010000000000",
		641 => "00000000000000000000000000000000",
		642 => "00000000000000000000000000000000",
		643 => "00000000000000000000000000000000",
		644 => "00000000000000000000000000000000",
		645 => "00000000000000000000000000000000",
		646 => "00000000000000000000000000000000",
		647 => "00000000000000000000000000000000",
		648 => "00000000000000000000000000000000",
		649 => "00000000000000000000000000000000",
		650 => "00000000000000000000000000000000",
		651 => "00000000000000000000000000000000",
		652 => "00000000000000000000000000000000",
		653 => "00000000000000000000000000000000",
		654 => "00000000000000000000000000000000",
		655 => "00000000000000000000000000000000",
		656 => "00000000000000000000000000000000",
		657 => "00000000000000000000000000000000",
		658 => "00000000000000000000000000000000",
		659 => "00000000000000000000000000000000",
		660 => "00000000000000000000000000000000",
		661 => "00000000000000000000000000000000",
		662 => "00000000000000000000000000000000",
		663 => "00000000000000000000000000000000",
		664 => "00000000000000000000000000000000",
		665 => "00000000000000000000000000000000",
		666 => "00000000000000000000000000000000",
		667 => "00000000000000000000000000000000",
		668 => "00000000000000000000000000000000",
		669 => "00000000000000000000000000000000",
		670 => "00000000000000000000000000000000",
		671 => "00000000000000000000000000000000",
		672 => "00000000000000000000000000000000",
		673 => "00000000000000000000000000000000",
		674 => "00000000000000000000000000000000",
		675 => "00000000000000000000000000000000",
		676 => "00000000000000000000000000000000",
		677 => "00000000000000000000000000000000",
		678 => "00000000000000000000000000000000",
		679 => "00000000000000000000000000000000",
		680 => "00000000000000000000000000000000",
		681 => "00000000000000000000000000000000",
		682 => "00000000000000000000000000000000",
		683 => "00000000000000000000000000000000",
		684 => "00000000000000000000000000000000",
		685 => "00000000000000000000000000000000",
		686 => "00000000000000000000000000000000",
		687 => "00000000000000000000000000000000",
		688 => "00000000000000000000000000000000",
		689 => "00000000000000000000000000000000",
		690 => "00000000000000000000000000000000",
		691 => "00000000000000000000000000000000",
		692 => "00000000000000000000000000000000",
		693 => "00000000000000000000000000000000",
		694 => "00000000000000000000000000000000",
		695 => "00000000000000000000000000000000",
		696 => "00000000000000000000000000000000",
		697 => "00000000000000000000000000000000",
		698 => "00000000000000000000000000000000",
		699 => "00000000000000000000000000000000",
		700 => "00000000000000000000000000000000",
		701 => "00000000000000000000000000000000",
		702 => "00000000000000000000000000000000",
		703 => "00000000000000000000000000000000",
		704 => "00000000000110000000010000000000",
		705 => "00000000000000000000000000000000",
		706 => "00000000000000000000000000000000",
		707 => "00000000000000000000000000000000",
		708 => "00000000000000000000000000000000",
		709 => "00000000000000000000000000000000",
		710 => "00000000000000000000000000000000",
		711 => "00000000000000000000000000000000",
		712 => "00000000000000000000000000000000",
		713 => "00000000000000000000000000000000",
		714 => "00000000000000000000000000000000",
		715 => "00000000000000000000000000000000",
		716 => "00000000000000000000000000000000",
		717 => "00000000000000000000000000000000",
		718 => "00000000000000000000000000000000",
		719 => "00000000000000000000000000000000",
		720 => "00000000000000000000000000000000",
		721 => "00000000000000000000000000000000",
		722 => "00000000000000000000000000000000",
		723 => "00000000000000000000000000000000",
		724 => "00000000000000000000000000000000",
		725 => "00000000000000000000000000000000",
		726 => "00000000000000000000000000000000",
		727 => "00000000000000000000000000000000",
		728 => "00000000000000000000000000000000",
		729 => "00000000000000000000000000000000",
		730 => "00000000000000000000000000000000",
		731 => "00000000000000000000000000000000",
		732 => "00000000000000000000000000000000",
		733 => "00000000000000000000000000000000",
		734 => "00000000000000000000000000000000",
		735 => "00000000000000000000000000000000",
		736 => "00000000000000000000000000000000",
		737 => "00000000000000000000000000000000",
		738 => "00000000000000000000000000000000",
		739 => "00000000000000000000000000000000",
		740 => "00000000000000000000000000000000",
		741 => "00000000000000000000000000000000",
		742 => "00000000000000000000000000000000",
		743 => "00000000000000000000000000000000",
		744 => "00000000000000000000000000000000",
		745 => "00000000000000000000000000000000",
		746 => "00000000000000000000000000000000",
		747 => "00000000000000000000000000000000",
		748 => "00000000000000000000000000000000",
		749 => "00000000000000000000000000000000",
		750 => "00000000000000000000000000000000",
		751 => "00000000000000000000000000000000",
		752 => "00000000000000000000000000000000",
		753 => "00000000000000000000000000000000",
		754 => "00000000000000000000000000000000",
		755 => "00000000000000000000000000000000",
		756 => "00000000000000000000000000000000",
		757 => "00000000000000000000000000000000",
		758 => "00000000000000000000000000000000",
		759 => "00000000000000000000000000000000",
		760 => "00000000000000000000000000000000",
		761 => "00000000000000000000000000000000",
		762 => "00000000000000000000000000000000",
		763 => "00000000000000000000000000000000",
		764 => "00000000000000000000000000000000",
		765 => "00000000000000000000000000000000",
		766 => "00000000000000000000000000000000",
		767 => "00000000000000000000000000000000",
		768 => "00000000000110000000010000000000",
		769 => "00000000000000000000000000000000",
		770 => "00000000000000000000000000000000",
		771 => "00000000000000000000000000000000",
		772 => "00000000000000000000000000000000",
		773 => "00000000000000000000000000000000",
		774 => "00000000000000000000000000000000",
		775 => "00000000000000000000000000000000",
		776 => "00000000000000000000000000000000",
		777 => "00000000000000000000000000000000",
		778 => "00000000000000000000000000000000",
		779 => "00000000000000000000000000000000",
		780 => "00000000000000000000000000000000",
		781 => "00000000000000000000000000000000",
		782 => "00000000000000000000000000000000",
		783 => "00000000000000000000000000000000",
		784 => "00000000000000000000000000000000",
		785 => "00000000000000000000000000000000",
		786 => "00000000000000000000000000000000",
		787 => "00000000000000000000000000000000",
		788 => "00000000000000000000000000000000",
		789 => "00000000000000000000000000000000",
		790 => "00000000000000000000000000000000",
		791 => "00000000000000000000000000000000",
		792 => "00000000000000000000000000000000",
		793 => "00000000000000000000000000000000",
		794 => "00000000000000000000000000000000",
		795 => "00000000000000000000000000000000",
		796 => "00000000000000000000000000000000",
		797 => "00000000000000000000000000000000",
		798 => "00000000000000000000000000000000",
		799 => "00000000000000000000000000000000",
		800 => "00000000000000000000000000000000",
		801 => "00000000000000000000000000000000",
		802 => "00000000000000000000000000000000",
		803 => "00000000000000000000000000000000",
		804 => "00000000000000000000000000000000",
		805 => "00000000000000000000000000000000",
		806 => "00000000000000000000000000000000",
		807 => "00000000000000000000000000000000",
		808 => "00000000000000000000000000000000",
		809 => "00000000000000000000000000000000",
		810 => "00000000000000000000000000000000",
		811 => "00000000000000000000000000000000",
		812 => "00000000000000000000000000000000",
		813 => "00000000000000000000000000000000",
		814 => "00000000000000000000000000000000",
		815 => "00000000000000000000000000000000",
		816 => "00000000000000000000000000000000",
		817 => "00000000000000000000000000000000",
		818 => "00000000000000000000000000000000",
		819 => "00000000000000000000000000000000",
		820 => "00000000000000000000000000000000",
		821 => "00000000000000000000000000000000",
		822 => "00000000000000000000000000000000",
		823 => "00000000000000000000000000000000",
		824 => "00000000000000000000000000000000",
		825 => "00000000000000000000000000000000",
		826 => "00000000000000000000000000000000",
		827 => "00000000000000000000000000000000",
		828 => "00000000000000000000000000000000",
		829 => "00000000000000000000000000000000",
		830 => "00000000000000000000000000000000",
		831 => "00000000000000000000000000000000",
		832 => "00000000000110000000010000000000",
		833 => "00000000000000000000000000000000",
		834 => "00000000000000000000000000000000",
		835 => "00000000000000000000000000000000",
		836 => "00000000000000000000000000000000",
		837 => "00000000000000000000000000000000",
		838 => "00000000000000000000000000000000",
		839 => "00000000000000000000000000000000",
		840 => "00000000000000000000000000000000",
		841 => "00000000000000000000000000000000",
		842 => "00000000000000000000000000000000",
		843 => "00000000000000000000000000000000",
		844 => "00000000000000000000000000000000",
		845 => "00000000000000000000000000000000",
		846 => "00000000000000000000000000000000",
		847 => "00000000000000000000000000000000",
		848 => "00000000000000000000000000000000",
		849 => "00000000000000000000000000000000",
		850 => "00000000000000000000000000000000",
		851 => "00000000000000000000000000000000",
		852 => "00000000000000000000000000000000",
		853 => "00000000000000000000000000000000",
		854 => "00000000000000000000000000000000",
		855 => "00000000000000000000000000000000",
		856 => "00000000000000000000000000000000",
		857 => "00000000000000000000000000000000",
		858 => "00000000000000000000000000000000",
		859 => "00000000000000000000000000000000",
		860 => "00000000000000000000000000000000",
		861 => "00000000000000000000000000000000",
		862 => "00000000000000000000000000000000",
		863 => "00000000000000000000000000000000",
		864 => "00000000000000000000000000000000",
		865 => "00000000000000000000000000000000",
		866 => "00000000000000000000000000000000",
		867 => "00000000000000000000000000000000",
		868 => "00000000000000000000000000000000",
		869 => "00000000000000000000000000000000",
		870 => "00000000000000000000000000000000",
		871 => "00000000000000000000000000000000",
		872 => "00000000000000000000000000000000",
		873 => "00000000000000000000000000000000",
		874 => "00000000000000000000000000000000",
		875 => "00000000000000000000000000000000",
		876 => "00000000000000000000000000000000",
		877 => "00000000000000000000000000000000",
		878 => "00000000000000000000000000000000",
		879 => "00000000000000000000000000000000",
		880 => "00000000000000000000000000000000",
		881 => "00000000000000000000000000000000",
		882 => "00000000000000000000000000000000",
		883 => "00000000000000000000000000000000",
		884 => "00000000000000000000000000000000",
		885 => "00000000000000000000000000000000",
		886 => "00000000000000000000000000000000",
		887 => "00000000000000000000000000000000",
		888 => "00000000000000000000000000000000",
		889 => "00000000000000000000000000000000",
		890 => "00000000000000000000000000000000",
		891 => "00000000000000000000000000000000",
		892 => "00000000000000000000000000000000",
		893 => "00000000000000000000000000000000",
		894 => "00000000000000000000000000000000",
		895 => "00000000000000000000000000000000",
		896 => "00000000000110000000010000000000",
		2048 => "11011000111000000100000000010010",
		2049 => "00111110001001110011100010001100",
		2050 => "11100000000010000000000000000000",
		2051 => "00001001000000001100000010001100",
		2052 => "11100000000001000000000000000000",
		2053 => "00001001110110001110000001000000",
		2054 => "00010010001111100010011100110001",
		2055 => "00111110001001110011100010001100",
		2056 => "11100000000010000000000000000000",
		2057 => "00001001010001111101001001001000",
		2058 => "00111000111000001000100000111110",
		2059 => "00100111001100001000110011000000",
		2060 => "00101000000000000000000000001001",
		2061 => "00111000110001100010000000111110",
		2062 => "00100111001100011101100011100000",
		2063 => "00000000000100100011111000100111",
		2064 => "00110000100011001100000000110000",
		2065 => "00000000000000000000100100000000",
		2066 => "11001111001111100010011100110001",
		2067 => "11001100110000000100110100000100",
		2068 => "00111110001001110011100010001100",
		2069 => "11100000001100000000000000000000",
		2070 => "00001001000001001110011010001100",
		2071 => "00000000000001000000000000000000",
		2072 => "00001001000011010100000010001100",
		2073 => "10100000000000000000000000000000",
		2074 => "00001001000000001111100000100100",
		2075 => "10100111000000000011111000000101",
		2076 => "00101001010000010000010101001111",
		2077 => "00000000111000001000110011100000",
		2078 => "00100000000000000000000000001001",
		2079 => "00000000111110001001110111000111",
		2080 => "01011001000000000000000000000000",
		2081 => "01000111001001001111111100000000",
		2082 => "11111111100011001110000000100000",
		2083 => "00000000000000000000100101000001",
		2084 => "00000111000111110000110101000000",
		2085 => "10001100111000000000000000000000",
		2086 => "00000000000010010000000011011000",
		2087 => "00100100111001100000000000111110",
		2088 => "00000111001110010100000100000111",
		2089 => "01001111000000001110100010001100",
		2090 => "11100000000011110000000000000000",
		
		2091 => "00001001000011000000000000000000", -- aqui � onde faz o byte enable mudar. original: 2091 => "00000000000010010000110000000000",

		
		
		2092 => "00000000000000000010000010110100",
		2093 => "01001000011001010110110001101100",
		2094 => "01101111001011000010000001010111",
		2095 => "01101111011100100110110001100100",
		2096 => "00100001000010100000000000000000",
		OTHERS => "00000000000000000000000000000000"
		-- OTHERS => (others=>'0') 
	);       
	


begin
    process(clk, addr)
    begin
	if( clk'event and clk = '1' ) then
		data_out <= dados(conv_integer(addr));
    end if;
    end process;
end Behav;

--------------------------------------------------------------