library verilog;
use verilog.vl_types.all;
entity ba22_top_qmem is
    port(
        clk_i           : in     vl_logic;
        rst_i           : in     vl_logic;
        iqmem_stb       : in     vl_logic;
        iqmem_we        : in     vl_logic;
        iqmem_addr      : in     vl_logic_vector(31 downto 0);
        iqmem_byte_en   : in     vl_logic_vector(3 downto 0);
        iqmem_wdata     : in     vl_logic_vector(31 downto 0);
        cpuid_i         : in     vl_logic_vector(31 downto 0);
        boot_devsel_i   : in     vl_logic;
        ben_le_sel_i    : in     vl_logic;
        dahb_clk_i      : in     vl_logic;
        dahb_rstn_i     : in     vl_logic;
        dahb_addr_o     : out    vl_logic_vector(31 downto 0);
        dahb_trans_o    : out    vl_logic_vector(1 downto 0);
        dahb_write_o    : out    vl_logic;
        dahb_size_o     : out    vl_logic_vector(2 downto 0);
        dahb_burst_o    : out    vl_logic_vector(2 downto 0);
        dahb_prot_o     : out    vl_logic_vector(3 downto 0);
        dahb_wdata_o    : out    vl_logic_vector(31 downto 0);
        dahb_rdata_i    : in     vl_logic_vector(31 downto 0);
        dahb_ready_i    : in     vl_logic;
        dahb_resp_i     : in     vl_logic_vector(1 downto 0);
        dahb_busreq_o   : out    vl_logic;
        dahb_lock_o     : out    vl_logic;
        dahb_grant_i    : in     vl_logic;
        dbg_stall_i     : in     vl_logic;
        dbg_ewt_i       : in     vl_logic;
        dbg_lss_o       : out    vl_logic_vector(3 downto 0);
        dbg_is_o        : out    vl_logic_vector(1 downto 0);
        dbg_wp_o        : out    vl_logic_vector(10 downto 0);
        dbg_bp_o        : out    vl_logic;
        dbg_stb_i       : in     vl_logic;
        dbg_we_i        : in     vl_logic;
        dbg_adr_i       : in     vl_logic_vector(15 downto 0);
        dbg_dat_i       : in     vl_logic_vector(31 downto 0);
        dbg_dat_o       : out    vl_logic_vector(31 downto 0);
        dbg_ack_o       : out    vl_logic;
        pic_int_i       : in     vl_logic_vector(2 downto 0);
        pm_clk_i        : in     vl_logic;
        pm_stall_i      : in     vl_logic;
        pm_stalled_o    : out    vl_logic;
        pm_clmode_i     : in     vl_logic_vector(7 downto 0);
        pm_event_o      : out    vl_logic;
        du_clk_i        : in     vl_logic;
        du_clk_en_o     : out    vl_logic;
        rf_clk_i        : in     vl_logic;
        rf_clk_en_o     : out    vl_logic
    );
end ba22_top_qmem;
