--------------------------------------------------------------
-- ROM - Template
-- Author: Renato Sampaio
-- Date: 21/02/2013
--------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;		 
use ieee.std_logic_unsigned.all;

entity ROM is
port(	clk   : in std_logic;
		addr	: in std_logic_vector(3 downto 0);
		data_out: out std_logic_vector(31 downto 0)
);
end ROM;

--------------------------------------------------------------

architecture Behav of ROM is

    type ROM_Array is array (0 to 2047) 
	of std_logic_vector(31 downto 0);

    constant dados: ROM_Array := (
		0 => "11111111110110101011110001110000",
		1 => "00000010001100011110011011010000",
		2 => "00000101000111111101100111010000",
		3 => "00001000110110101111110100000000",
		4 => "00001101000001100100110011000000",
		5 => "00010001110001110100101111110000",
		6 => "00010110001111111101110100110000",
		7 => "00011010100111110110110011100000",
		8 => "00011111011111100101000011100000",
		9 => "00100100110001111010111111000000",
		10 => "00101010101011110000101001010000",
		11 => "00110001001010000011000010110000",
		12 => "00110111101001010110000110100000",
		13 => "00111100110000101011010100010000",
		14 => "01000000100101100111001000110000",
		15 => "01000011010101111011001101010000",
		OTHERS => "00000000000000000000000000000000"
	);       

begin
    process(clk, addr)
    begin
	if( clk'event and clk = '1' ) then
		data_out <= dados(conv_integer(addr));
    end if;
    end process;
end Behav;

--------------------------------------------------------------